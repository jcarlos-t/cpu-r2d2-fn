`timescale 1ns / 1ps

module testbench_matmul();
  // Señales del DUT (Device Under Test)
  logic        clk;
  logic        reset;
  logic [31:0] WriteDataM, DataAdrM;
  logic        MemWriteM;
  
  logic [31:0] PCF;
  logic [31:0] InstrF;
  logic [31:0] pc_backup;
  logic        save_pc;
  logic        save_pc;
  logic        im_sel;
  logic        toggle_fsm;
  logic        fsm_state;
  
  // Variables para control de test
  integer cycle_count;
  
  // Instancia del DUT
  top dut(
    .clk(clk),
    .reset(reset),
    .WriteDataM(WriteDataM),
    .DataAdrM(DataAdrM),
    .MemWriteM(MemWriteM),
    .file_name("program.mem")  // Archivo de programa principal
  );
  
  // Generación de reloj: 10ns periodo (100MHz)
  initial begin
    clk = 0;
    forever #5 clk = ~clk;
  end
  
  // Asignación de señales internas mediante hierarchical reference
  assign PCF = dut.PCF;
  assign InstrF = dut.InstrF;
  
  // Señales de MATMUL - ahora con las rutas correctas
  assign pc_backup = dut.pc_backup;
  assign save_pc = dut.save_pc;
  assign im_sel = dut.im_sel;
  assign toggle_fsm = dut.toggle_fsm;
  assign fsm_state = dut.fsm.state;
  
  // Secuencia de reset y test
  initial begin
    $display("================================================================================");
    $display("  TESTBENCH MATMUL - Verificación de Microcodigo");
    $display("================================================================================");
    $display("\n[HEADER] Señales principales de control:");
    $display("  FSM_STATE: Estado actual del FSM (0=NORMAL, 1=MATMUL2)");
    $display("  IM_SEL: Selección de instruction memory (0=normal, 1=matmul2)");
    $display("  SAVE_PC: Habilita guardado de PC");
    $display("  RESET_PC: Resetea PC a 0");
    $display("================================================================================\n");
    
    // Inicialización
    cycle_count = 0;
    reset = 1;
    
    // Mantener reset por 2 ciclos
    #20;
    reset = 0;
    
    $display("[INFO] Reset liberado, iniciando ejecución...\n");
    
    // Ejecutar por 200 ciclos de reloj
    repeat(200) begin
      @(posedge clk);
      cycle_count = cycle_count + 1;
    end
    
    $display("\n================================================================================");
    $display("  Test completado después de %0d ciclos", cycle_count);
    $display("================================================================================");
    $finish;
  end
  
  // Monitor detallado de señales en cada ciclo
  always @(posedge clk) begin
    if (!reset) begin
      $display("[CICLO %3d] PC=%08h | Instr=%08h | FSM=%b | IM_SEL=%b | WB: RegWr=%b Rd=%2d Val=%08h",
               cycle_count, PCF, InstrF, fsm_state, im_sel, 
               dut.riscv.RegWriteW, dut.riscv.RdW, dut.riscv.ResultW);
      
      // Monitor adicional para debug de datos
      if (fsm_state == 1'b1) begin
         $display("    [DEBUG] FP ALU: A=%h B=%h -> Res=%h", 
                  dut.riscv.dp.SrcAE_fp, dut.riscv.dp.SrcBE_fp, dut.riscv.dp.fpuResult);
         $display("    [DEBUG] Shadow Regs: x30(A)=%h, x31(B)=%h, x29(C)=%h",
                  dut.riscv.rf_int.rf[30], dut.riscv.rf_int.rf[31], dut.riscv.rf_int.rf[29]);
      end
    end
  end
  
  
  // Monitor de señales de control MATMUL con estado detallado
  always @(posedge clk) begin
    if (!reset) begin
      // Detectar inicio de MATMUL (Toggle en estado NORMAL)
      if (toggle_fsm && fsm_state == 1'b0) begin
        $display("\n╔═══════════════════════════════════════════════════════════════════╗");
        $display("║ >>> [MATMUL START] Ciclo %0d: STARTMATMUL2 detectado", 
                 cycle_count);
        $display("║     PC actual guardado: %08h", PCF);
        $display("║     PC+4 a guardar: %08h", PCF + 4);
        $display("║     Control: save_pc=%b, im_sel=%b, toggle_fsm=%b", 
                 save_pc, im_sel, toggle_fsm);
        $display("║     FSM: Estado actual=%b, próximo estado=MATMUL2(1)",
                 fsm_state);
        $display("╚═══════════════════════════════════════════════════════════════════╝\n");
      end
      
      // Detectar fin de MATMUL (Toggle en estado MATMUL2)
      if (toggle_fsm && fsm_state == 1'b1) begin
        $display("\n╔═══════════════════════════════════════════════════════════════════╗");
        $display("║ <<< [MATMUL END] Ciclo %0d: ENDMATMUL detectado", cycle_count);
        $display("║     Estado FSM actual: %b (%s)", fsm_state,
                 fsm_state == 1'b1 ? "MATMUL2" : "NORMAL");
        $display("║     PC backup a restaurar: %08h", pc_backup);
        $display("║     Retornando a flujo normal...");
        $display("╚═══════════════════════════════════════════════════════════════════╝\n");
      end
    end
  end
  
  
  // Monitor de escrituras a memoria
  always @(posedge clk) begin
    if (!reset && MemWriteM) begin
      $display("\n    [MEM WRITE] Dirección: %08h, Dato: %08h (Ciclo %0d)",
               DataAdrM, WriteDataM, cycle_count);
    end
  end
  
  // Monitor de cambios en el PC
  logic [31:0] prev_pc;
  initial prev_pc = 0;
  
  always @(posedge clk) begin
    if (!reset) begin
      if (PCF != prev_pc + 4 && cycle_count > 0) begin
        $display("\n    [PC JUMP] De %08h a %08h (diferencia: %0d) en ciclo %0d",
                 prev_pc, PCF, $signed(PCF - prev_pc), cycle_count);
      end
      prev_pc = PCF;
    end
  end
  
  // Generación de archivo VCD para GTKWave (opcional)
  initial begin
    $dumpfile("testbench_matmul.vcd");
    $dumpvars(0, testbench_matmul);
    $dumpvars(0, dut);
  end
  
  // Monitor de instrucciones decodificadas
  logic [6:0] opcode;
  assign opcode = InstrF[6:0];
  
  always @(posedge clk) begin
    if (!reset && cycle_count > 0) begin
      case (opcode)
        7'b1111010: begin
          if (InstrF[14:12] == 3'b000) $display("\n>>> [DECODE] STARTMATMUL2 detectado en ciclo %0d", cycle_count);
          else if (InstrF[14:12] == 3'b111) $display("\n<<< [DECODE] ENDMATMUL detectado en ciclo %0d", cycle_count);
        end
        7'b0110011: if (cycle_count % 10 == 0) $display("    [DECODE] R-type (Integer)");
        7'b1010011: if (cycle_count % 10 == 0) $display("    [DECODE] R-type (FPU)");
        7'b0000011: if (cycle_count % 10 == 0) $display("    [DECODE] LW");
        7'b0100011: if (cycle_count % 10 == 0) $display("    [DECODE] SW");
        7'b1100011: if (cycle_count % 10 == 0) $display("    [DECODE] BEQ");
        7'b1101111: $display("    [DECODE] JAL en ciclo %0d", cycle_count);
      endcase
    end
  end
  
  // Timeout de seguridad
  initial begin
    #100000; // 100us timeout
    $display("\n[ERROR] TIMEOUT - El test excedió el tiempo máximo de ejecución");
    $finish;
  end

endmodule
